RC discharge circuit
R1 0 1 100
C1 1 0 10u IC=10
.TRAN 1E-6 5E-3