PWL source and resistor circuit
V1 1 0 PWL(0.5u 2 2u -1 5u 0 9u 7)
R1 0 1 100
.TRAN 1n 10u