Sine source and resistor circuit
V1 1 0 SIN(0 1 60 0.002083333)
R1 0 1 100
.TRAN 1E-5 5E-2