RC discharge circuit
R1 0 1 100
L1 1 0 10u IC=0.1
.TRAN 1E-10 5E-7